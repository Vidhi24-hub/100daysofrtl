//Clock Generator having 10MHz frequency
'timescale 10ns/10ps

module clk_gen(clk);
  input clk;
endmodule